module cpu_datapath
(

);



endmodule
