module lda_control
(
  input clk,
  input reset,
  
  input i_start,
  
  output o_done,
  
  output o_plot,
  
  input i_x0_gt_x1,
  
  output o_ld_constants,
  output o_ld_error,
  output o_ld_ystep,
  output o_ld_xstep,
  output o_ld_y,
  output o_ld_x
);



endmodule
