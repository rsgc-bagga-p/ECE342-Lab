module lda_control
(


);



endmodule
