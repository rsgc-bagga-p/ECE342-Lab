module lda_asc_datapath
(
  input i_clk,
  input i_reset


);



endmodule
