module alu
(

);



endmodule
