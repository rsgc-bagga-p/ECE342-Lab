module lda_datapath
(


);



endmodule
