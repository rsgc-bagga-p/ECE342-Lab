module led_ctrl
(
	input clk,
	input reset,

	input i_val,
	input i_enable,
	output logic o_out
);

	always_ff @ (posedge clk or posedge reset) begin
		if (reset) o_out <= '0;
		else if (i_enable) o_out <= i_val;
	end

endmodule
