module cpu_control
(
  input i_clk,
  input i_reset
);



endmodule
