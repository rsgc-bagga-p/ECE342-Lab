`timescale 100ps/100ps // Makes 50GHz

module tb_asc();



endmodule
