module cpu_control
(

);



endmodule
